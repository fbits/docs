[{"type":"Conceptual","source_relative_path":"articles/intro.md","output":{".html":{"relative_path":"articles/intro.html","link_to_path":"/github/workspace/docfx_project/obj/.cache/build/ii5uv0ri.izo/733w16kd.zwp","hash":"oulplDd4bW8jlLrrtORwAQ=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"index.md","output":{".html":{"relative_path":"index.html","link_to_path":"/github/workspace/docfx_project/obj/.cache/build/ii5uv0ri.izo/7uemy0ft.cyw","hash":"SkaVYJvbwK6YgkAXK4s2ow=="}},"is_incremental":true,"version":""},{"type":"Conceptual","source_relative_path":"api/index.md","output":{".html":{"relative_path":"api/index.html","link_to_path":"/github/workspace/docfx_project/obj/.cache/build/ii5uv0ri.izo/jamla758.nqq","hash":"EFBUNp8nfORMMT/9qfaDXg=="}},"is_incremental":true,"version":""},{"type":"Toc","source_relative_path":"articles/toc.yml","output":{".html":{"relative_path":"articles/toc.html","link_to_path":"/github/workspace/docfx_project/obj/.cache/build/ii5uv0ri.izo/stgdq84p.td8","hash":"t7iiFrmuYmrKWisdq+lN6Q=="}},"is_incremental":false,"version":""},{"type":"Toc","source_relative_path":"toc.yml","output":{".html":{"relative_path":"toc.html","link_to_path":"/github/workspace/docfx_project/obj/.cache/build/ii5uv0ri.izo/0r5aheit.nta","hash":"k+/dkjFuwAVS32HduMpmBw=="}},"is_incremental":false,"version":""},{"type":"Toc","source_relative_path":"api/toc.yml","output":{".html":{"relative_path":"api/toc.html","link_to_path":"/github/workspace/docfx_project/obj/.cache/build/ii5uv0ri.izo/0fft5kk4.2io","hash":"eWl/m2iB2mgjZPbLc4xDqw=="}},"is_incremental":false,"version":""}]